** Profile: "SCHEMATIC1-vdc"  [ E:\An2_Sem2\Tehnici_CAD\Proiect\main-pspicefiles\schematic1\vdc.sim ] 

** Creating circuit file "vdc.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dimesionare_led.lib" 
.LIB "../../../main-pspicefiles/main.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM SET 0 1 0.05 
.WCASE DC v([OUT]) YMAX VARY BOTH  HI 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
