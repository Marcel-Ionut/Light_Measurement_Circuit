** Profile: "SCHEMATIC1-vac"  [ E:\An2_Sem2\Tehnici_CAD\Proiect\main-pspicefiles\schematic1\vac.sim ] 

** Creating circuit file "vac.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dimesionare_led.lib" 
.LIB "../../../main-pspicefiles/main.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 
.MC 10 TRAN v([OUT]) YMAX OUTPUT RUNS  SEED=200 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
